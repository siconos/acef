LINEAR_DC_CKT.CIR - SIMPLE CIRCUIT FOR NODAL ANALYSIS
*
VS	0	1	AC      1       SIN(0   1       1000)

*
R1	1	2	100
C1	2	3	0.02
L1	3	0	0.03
*
* ANALYSIS
.TRAN 	0.1us  10000uS
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(3)
.PROBE
.END
