RLMOS.CIR - SIMPLE CIRCUIT MOS test
*
*VIN	1	0	AC	1	SIN(0	10	2)
VIN1	1	0	DC	1
VIN2	2	0	DC	10

.model nmos nmos level=1 tox=100e-09 vto=2.0 kp=10.0
M1	2	1	3	0	nmos	w=0.0001	l=0.0001
R1	3 4 1
L1	4	0	0.0001
R2	4 0 1
*
.ic V(2)=10
.ic V(1)=1


*
* ANALYSIS
.TRAN 	0.01S  1S
* VIEW RESULTS
.PRINT	TRAN 	 V(3,4) V(1)	V(2)	V(3) V(4)
.PROBE
.END
