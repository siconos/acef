LINEAR_DC_CKT.CIR - SIMPLE CIRCUIT FOR NODAL ANALYSIS
*
VS	0	1	DC	2
IS	0	1	DC	1
*
R1	0	1	1000
C1	0	1	0.001
L1	1	0	0.002
*
* ANALYSIS
.TRAN 	1MS  10MS
* VIEW RESULTS
.PRINT	TRAN 	V(1)
.PROBE
.END
