BuckConverterRegul2


ValimI 1 0 3

* power mosfets : no cross conduction thanks to sum of Vt 
.model nmos nmos level=1 tox=100e-09 vto=2.0 kp=10.0
.model pmos pmos level=1 tox=100e-09 vto=-2.0 kp=10.0
mosnswitch 2 7 0 0 nmos w=0.0001 l=0.0001
mospswitch 2 7 1 1 pmos w=0.0001 l=0.0001


L1 2 3 10u
C1 3 0 22u
Rload 3 0 10.0

*Vbruit 33 0 PULSE(0 -1.8 0.1e-3 0.1e-4 0.1e-4 5e-9 )
*Vramp 6 0 PULSE(0 2.25 0 1.660e-6 5e-9 1e-9 1.6667e-6)

* these values of L1,C1 give a sliding mode
* L1 2 3 4u
* C1 3 0 10u

.MODEL DIODEDEF D N=1

Dnswitch 0 2 DIODEDEF
Dpswitch 2 1 DIODEDEF

Vramp 6 0 PULSE(0 2.25 0 1.660e-6 5e-9 1e-9 1.6667e-6)
*Vramp 6 0 PULSE(0 2.25 0 3e-6 5e-9 1e-9 3e-6)

Vref 4 0 PULSE(0 1.8 0 1e-4)

* first set of compensator parameters R11 R21 C11
R11 3 12 15.58E3
R21 13 11 5.613E6
C11 12 11 20E-12

* second set of compensator parameters R11 R21 C11
* R11 3 12 10E3
* R21 13 11 8E6
* C11 12 11 10E-12

R12 3 11 227.8E3
C21 5 13 1.9E-12

* amplifier
Eampli 14 0 4 11 10000.0
Ramp 14 5 1
Camp 5 0 5.305E-9

* comparator
*Bcomp 7 0 V=1.5*(tanh(10.0*V(6,5)) + 1.0)
.comp 6 5 7 Vmin=0 Vmax=3 Vepsilon=0.15

.options method=trap RELTOL=0.04

.save  v(3) v(2) 

.tran 50ps 0.0002
*.tran 50ps 50000000ps
.print tran  v(1) v(2) v(3) v(4) v(5) v(6) v(7) v(9) v(10) v(11) v(12) v(13) v(14) v(3,2)

.control
set width = 230
set nobreak
rusage everything
.endc
.end
