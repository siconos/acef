diode bridge

.subckt resis n1 n2
RresisName n1 n2 1000
.ends

C1 1 0 1uF
L1 1 0 10mH

xR1 2 3 resis

.MODEL DIODEDEF D N=0.25
DF1 1 2 DIODEDEF 
DR2 3 1 DIODEDEF 
DR1 0 2 DIODEDEF 
DF2 3 0 DIODEDEF 

.ic V(1)=10
.ic V(2)=10

.options method=trap RELTOL=0.04

.save  v(2)-V(3)

#.tran 1e-9 3e-4
.tran 1e-6 5e-3
.print tran 	v(2,3)

.control
set width = 230
set nobreak
rusage everything
.endc
.end
