LINEAR_DC_CKT.CIR - SIMPLE CIRCUIT FOR NODAL ANALYSIS
*
IS	0	1	DC	1A
*
C1	1	0	0.01
L1	1	0	0.02
*
* ANALYSIS
.TRAN 	1MS  10MS
* VIEW RESULTS
.PRINT	TRAN 	V(1)
.PROBE
.END
