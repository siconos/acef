RMOS.CIR - SIMPLE CIRCUIT MOS test
*
VIN	1	0	AC	1	SIN(0	3	2)
R1	2	0	10
V2	3	0	DC	1
*

.model nmos nmos level=1 tox=100e-09 vto=2.0 kp=10.0
M1	2	1	3	0	nmos	w=0.0001	l=0.0001

*
* ANALYSIS
.TRAN 	0.01S  1S
* VIEW RESULTS
.PRINT	TRAN 	V(1)	V(2)	V(3)
.PROBE
.END
