diode bridge

C1 1 0 1uF
L1 1 0 10mH
R1 2 3 1000

.MODEL DIODEDEF D N=0.25
DF1 1 2 DIODEDEF 
DR2 3 1 DIODEDEF 
DR1 0 2 DIODEDEF 
DF2 3 0 DIODEDEF 

.ic V(1)=10
.options method=trapezoidal

.control
set width = 140
set nobreak

tran 100u 10.0m uic
print col v(1) v(3) v(2,3) v(2) 
.endc

.END
