LINEAR_DC_CKT.CIR - SIMPLE CIRCUIT FOR NODAL ANALYSIS
*
VS	0	1	AC      1       SIN(0   1       1000)
*
R2	1	2	100
C1	2	0	2u
*
* ANALYSIS
.TRAN 	0.1us  10000uS
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2)
.PROBE
.END
