
*                                  3
*                           /--R1--.--->|------
* 5        1         2     /
* |----||---.---L----.----/
* |                       \
* |                        \
* |                         \
* VS                         |
* |                          |
* |                          R2
* |                          |
* |                          |
* |                         4.
* |                          |
* |                          |
* |                          |
* |                          \/
* |                          --
* |                          |
* |                          |
*
*
*

L1 1 2 10mH
R1 2 3 1000
R2 2 4 500

C1 1 5 1uF
VS	0	5	AC      1       SIN(0   1       1000)

.MODEL DIODEDEF D N=0.25
D1 3 0 DIODEDEF 
D2 0 4 DIODEDEF 

*.ic V(1)=10



* ANALYSIS
.TRAN 	0.1us  5000uS
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(3) V(4) V(5)
.PROBE
.END

